//test hello world for verilog  
module hello;
  initial
    begin
      $display("Hello, World");
      $finish ;
    end

    